library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY PGCD IS
PORT 
( 
	CLK      : in  STD_LOGIC;
	RESET    : in  STD_LOGIC;

	idata_a  : in  STD_LOGIC_VECTOR (31 downto 0);
	idata_b  : in  STD_LOGIC_VECTOR (31 downto 0);
	idata_en : in  STD_LOGIC;

	odata    : out STD_LOGIC_VECTOR (31 downto 0);
	odata_en : out STD_LOGIC
);
END PGCD;

architecture Behavioral of PGCD is
    TYPE STATE_TYPE IS (init, compute, output);
    SIGNAL current_state, next_state : STATE_TYPE;
    
    signal A     : signed(31 downto 0);
    signal B     : signed(31 downto 0);
    signal A1    : signed(31 downto 0);
    signal B1    : signed(31 downto 0);
    signal cpt   : unsigned(7 downto 0);

begin
    --State register
    PROCESS (CLK, RESET)
    BEGIN
        IF RESET = '1' THEN
            current_state  <= init;
        ELSIF (CLK'EVENT AND CLK = '1') THEN
            current_state <= next_state;
        END IF;
    END PROCESS;

    --next state
    PROCESS(current_state, A, B)
    begin
        case current_state is
            when init => 
                if (idata_en = '1') THEN
                    --inputs asserts
                    assert (A >= 0) report "idata_a < 0" severity failure;
                    assert (B >= 0) report "idata_b < 0" severity failure;
                    assert (A <= 65535) report "idata_a > 65535" severity failure;
                    assert (B <= 65535) report "idata_b > 65535" severity failure;
                    
                    A1 <= signed(idata_a);
                    B1 <= signed(idata_b);
                    next_state <= compute;
                else 
                    next_state <= current_state;
                end if;
                
            when compute =>
                assert (idata_en = '0') report "Load while computing" severity failure;
                
                if (A = B) then
                    next_state <= output;
                else
                    next_state <= current_state;
                end if;
                    
            when output => 
                --pragma translate_off
                REPORT "cpt = " & integer'image(to_integer( cpt ));
                --pragma translate_on

                --outputs asserts
                assert (idata_en = '0') report "Load while getting outputs" severity failure;
                assert (A1 >= A) report "Output bigger than input" severity failure;
                assert (B1 >= B) report "Output bigger than input" severity failure;
                assert (A >= 0) report "Negative output" severity failure;
                next_state <= init;
        end case;
    end process;

    --output
    process(current_state, A)
    begin
        case current_state is
            when init | compute =>  odata_en    <= '0';
                                    odata       <= std_logic_vector(A);
                        
            when output =>          odata_en    <= '1';
                                    odata       <= std_logic_vector(A);
        end case;
    end process;

    --compute pgcd
    process(CLK, RESET, current_state)
    begin
        IF (RESET = '1') THEN
            A   <= (others => '0');
            B   <= (others => '0');
            A1  <= (others => '0');
            B1  <= (others => '0');

        elsif (current_state = init) then
            A  <= signed(idata_a);
            B  <= signed(idata_b);
            A1 <= signed(idata_a);
            B1 <= signed(idata_b);
            cpt <= to_unsigned(0, cpt'length);

        ELSIF (CLK'EVENT AND CLK = '1' AND current_state = compute) THEN
            cpt <= cpt + 1;

            if (A = 0) then
                A <= B;
            elsif (B = 0) then
                B <= A;
            
            elsif (A > (B(27 downto 0) & "0000")) then
                A <= A - (B(27 downto 0) & "0000");
            elsif (B > (A(27 downto 0) & "0000")) then
                B <= B - (A(27 downto 0) & "0000");
            
            elsif (A > B) then 
                A <= A - B;
            elsif (B > A) then 
                B <= B - A;
            end if;
        end if;
    end process;

end Behavioral;